-------------------------------------------------------------------------------
-- Dr. Kaputa & Adam Hemmouda
-- single bit full adder test bench
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;      -- gives you the std_logic type

entity full_adder_single_bit_str_tb is 
end full_adder_single_bit_str_tb;

architecture arch of full_adder_single_bit_str_tb is

component full_adder_single_bit_str
  port(
    a      : in std_logic;    -- Input (A)
    b      : in std_logic;    -- Input (B)
    cin     : in std_logic;   -- Input (CIN)
    sum     : out std_logic;  -- Output (SUM)
    cout    : out std_logic   -- Output (COUT)
    );
  end component;
  
signal a    : std_logic := '0';
signal b    : std_logic := '0'; 
signal cin  : std_logic := '0';
signal sum  : std_logic;
signal cout : std_logic;

begin 
  uut: full_adder_single_bit_str 
    port map(
      a     => a,
      b     => b,
      cin   => cin,
      sum   => sum,
      cout  => cout
    );

  a <= not a after 10 ns;
  b <= not b after 20 ns;
  cin <= not cin after 40 ns;
end arch;